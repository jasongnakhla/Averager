----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 11/10/2020 12:34:46 AM
-- Design Name: 
-- Module Name: DWPP - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity DWPP is
    Port ( clk : in STD_LOGIC;
           rst: in STD_LOGIC;
           d : in STD_LOGIC_VECTOR(8 downto 0);
           q_hadder : out STD_LOGIC_VECTOR(7 downto 0);
           q_product : out STD_LOGIC_VECTOR(15 downto 0));
end DWPP;

architecture Behavioral of DWPP is

signal temp: STD_LOGIC_VECTOR(16 downto 0):=(others=>'0');

begin
process(clk,rst,d)
    begin
    if (rst='1') then
        temp <= (others => '0');
    elsif(rising_edge(clk)) then
        temp <= d & temp(9 downto 2);
    end if;
end process;

q_hadder <= '0' & temp(16 downto 10); 
q_product <= temp(15 downto 0); 

end Behavioral;

